module Float_8bit_Table(U, F, P);
	input [7:0] U;
	output reg [7:0] F;
	output reg [2:0] P;
	
	reg [10:0] Table[0:255];
	
	initial begin
		Table[0]=11'b00000000000;
		Table[1]=11'b10000000000;
		Table[2]=11'b10000000001;
		Table[3]=11'b11000000001;
		Table[4]=11'b10000000010;
		Table[5]=11'b10100000010;
		Table[6]=11'b11000000010;
		Table[7]=11'b11100000010;
		Table[8]=11'b10000000011;
		Table[9]=11'b10010000011;
		Table[10]=11'b10100000011;
		Table[11]=11'b10110000011;
		Table[12]=11'b11000000011;
		Table[13]=11'b11010000011;
		Table[14]=11'b11100000011;
		Table[15]=11'b11110000011;
		Table[16]=11'b10000000100;
		Table[17]=11'b10001000100;
		Table[18]=11'b10010000100;
		Table[19]=11'b10011000100;
		Table[20]=11'b10100000100;
		Table[21]=11'b10101000100;
		Table[22]=11'b10110000100;
		Table[23]=11'b10111000100;
		Table[24]=11'b11000000100;
		Table[25]=11'b11001000100;
		Table[26]=11'b11010000100;
		Table[27]=11'b11011000100;
		Table[28]=11'b11100000100;
		Table[29]=11'b11101000100;
		Table[30]=11'b11110000100;
		Table[31]=11'b11111000100;
		Table[32]=11'b10000000101;
		Table[33]=11'b10000100101;
		Table[34]=11'b10001000101;
		Table[35]=11'b10001100101;
		Table[36]=11'b10010000101;
		Table[37]=11'b10010100101;
		Table[38]=11'b10011000101;
		Table[39]=11'b10011100101;
		Table[40]=11'b10100000101;
		Table[41]=11'b10100100101;
		Table[42]=11'b10101000101;
		Table[43]=11'b10101100101;
		Table[44]=11'b10110000101;
		Table[45]=11'b10110100101;
		Table[46]=11'b10111000101;
		Table[47]=11'b10111100101;
		Table[48]=11'b11000000101;
		Table[49]=11'b11000100101;
		Table[50]=11'b11001000101;
		Table[51]=11'b11001100101;
		Table[52]=11'b11010000101;
		Table[53]=11'b11010100101;
		Table[54]=11'b11011000101;
		Table[55]=11'b11011100101;
		Table[56]=11'b11100000101;
		Table[57]=11'b11100100101;
		Table[58]=11'b11101000101;
		Table[59]=11'b11101100101;
		Table[60]=11'b11110000101;
		Table[61]=11'b11110100101;
		Table[62]=11'b11111000101;
		Table[63]=11'b11111100101;
		Table[64]=11'b10000000110;
		Table[65]=11'b10000010110;
		Table[66]=11'b10000100110;
		Table[67]=11'b10000110110;
		Table[68]=11'b10001000110;
		Table[69]=11'b10001010110;
		Table[70]=11'b10001100110;
		Table[71]=11'b10001110110;
		Table[72]=11'b10010000110;
		Table[73]=11'b10010010110;
		Table[74]=11'b10010100110;
		Table[75]=11'b10010110110;
		Table[76]=11'b10011000110;
		Table[77]=11'b10011010110;
		Table[78]=11'b10011100110;
		Table[79]=11'b10011110110;
		Table[80]=11'b10100000110;
		Table[81]=11'b10100010110;
		Table[82]=11'b10100100110;
		Table[83]=11'b10100110110;
		Table[84]=11'b10101000110;
		Table[85]=11'b10101010110;
		Table[86]=11'b10101100110;
		Table[87]=11'b10101110110;
		Table[88]=11'b10110000110;
		Table[89]=11'b10110010110;
		Table[90]=11'b10110100110;
		Table[91]=11'b10110110110;
		Table[92]=11'b10111000110;
		Table[93]=11'b10111010110;
		Table[94]=11'b10111100110;
		Table[95]=11'b10111110110;
		Table[96]=11'b11000000110;
		Table[97]=11'b11000010110;
		Table[98]=11'b11000100110;
		Table[99]=11'b11000110110;
		Table[100]=11'b11001000110;
		Table[101]=11'b11001010110;
		Table[102]=11'b11001100110;
		Table[103]=11'b11001110110;
		Table[104]=11'b11010000110;
		Table[105]=11'b11010010110;
		Table[106]=11'b11010100110;
		Table[107]=11'b11010110110;
		Table[108]=11'b11011000110;
		Table[109]=11'b11011010110;
		Table[110]=11'b11011100110;
		Table[111]=11'b11011110110;
		Table[112]=11'b11100000110;
		Table[113]=11'b11100010110;
		Table[114]=11'b11100100110;
		Table[115]=11'b11100110110;
		Table[116]=11'b11101000110;
		Table[117]=11'b11101010110;
		Table[118]=11'b11101100110;
		Table[119]=11'b11101110110;
		Table[120]=11'b11110000110;
		Table[121]=11'b11110010110;
		Table[122]=11'b11110100110;
		Table[123]=11'b11110110110;
		Table[124]=11'b11111000110;
		Table[125]=11'b11111010110;
		Table[126]=11'b11111100110;
		Table[127]=11'b11111110110;
		Table[128]=11'b10000000111;
		Table[129]=11'b10000001111;
		Table[130]=11'b10000010111;
		Table[131]=11'b10000011111;
		Table[132]=11'b10000100111;
		Table[133]=11'b10000101111;
		Table[134]=11'b10000110111;
		Table[135]=11'b10000111111;
		Table[136]=11'b10001000111;
		Table[137]=11'b10001001111;
		Table[138]=11'b10001010111;
		Table[139]=11'b10001011111;
		Table[140]=11'b10001100111;
		Table[141]=11'b10001101111;
		Table[142]=11'b10001110111;
		Table[143]=11'b10001111111;
		Table[144]=11'b10010000111;
		Table[145]=11'b10010001111;
		Table[146]=11'b10010010111;
		Table[147]=11'b10010011111;
		Table[148]=11'b10010100111;
		Table[149]=11'b10010101111;
		Table[150]=11'b10010110111;
		Table[151]=11'b10010111111;
		Table[152]=11'b10011000111;
		Table[153]=11'b10011001111;
		Table[154]=11'b10011010111;
		Table[155]=11'b10011011111;
		Table[156]=11'b10011100111;
		Table[157]=11'b10011101111;
		Table[158]=11'b10011110111;
		Table[159]=11'b10011111111;
		Table[160]=11'b10100000111;
		Table[161]=11'b10100001111;
		Table[162]=11'b10100010111;
		Table[163]=11'b10100011111;
		Table[164]=11'b10100100111;
		Table[165]=11'b10100101111;
		Table[166]=11'b10100110111;
		Table[167]=11'b10100111111;
		Table[168]=11'b10101000111;
		Table[169]=11'b10101001111;
		Table[170]=11'b10101010111;
		Table[171]=11'b10101011111;
		Table[172]=11'b10101100111;
		Table[173]=11'b10101101111;
		Table[174]=11'b10101110111;
		Table[175]=11'b10101111111;
		Table[176]=11'b10110000111;
		Table[177]=11'b10110001111;
		Table[178]=11'b10110010111;
		Table[179]=11'b10110011111;
		Table[180]=11'b10110100111;
		Table[181]=11'b10110101111;
		Table[182]=11'b10110110111;
		Table[183]=11'b10110111111;
		Table[184]=11'b10111000111;
		Table[185]=11'b10111001111;
		Table[186]=11'b10111010111;
		Table[187]=11'b10111011111;
		Table[188]=11'b10111100111;
		Table[189]=11'b10111101111;
		Table[190]=11'b10111110111;
		Table[191]=11'b10111111111;
		Table[192]=11'b11000000111;
		Table[193]=11'b11000001111;
		Table[194]=11'b11000010111;
		Table[195]=11'b11000011111;
		Table[196]=11'b11000100111;
		Table[197]=11'b11000101111;
		Table[198]=11'b11000110111;
		Table[199]=11'b11000111111;
		Table[200]=11'b11001000111;
		Table[201]=11'b11001001111;
		Table[202]=11'b11001010111;
		Table[203]=11'b11001011111;
		Table[204]=11'b11001100111;
		Table[205]=11'b11001101111;
		Table[206]=11'b11001110111;
		Table[207]=11'b11001111111;
		Table[208]=11'b11010000111;
		Table[209]=11'b11010001111;
		Table[210]=11'b11010010111;
		Table[211]=11'b11010011111;
		Table[212]=11'b11010100111;
		Table[213]=11'b11010101111;
		Table[214]=11'b11010110111;
		Table[215]=11'b11010111111;
		Table[216]=11'b11011000111;
		Table[217]=11'b11011001111;
		Table[218]=11'b11011010111;
		Table[219]=11'b11011011111;
		Table[220]=11'b11011100111;
		Table[221]=11'b11011101111;
		Table[222]=11'b11011110111;
		Table[223]=11'b11011111111;
		Table[224]=11'b11100000111;
		Table[225]=11'b11100001111;
		Table[226]=11'b11100010111;
		Table[227]=11'b11100011111;
		Table[228]=11'b11100100111;
		Table[229]=11'b11100101111;
		Table[230]=11'b11100110111;
		Table[231]=11'b11100111111;
		Table[232]=11'b11101000111;
		Table[233]=11'b11101001111;
		Table[234]=11'b11101010111;
		Table[235]=11'b11101011111;
		Table[236]=11'b11101100111;
		Table[237]=11'b11101101111;
		Table[238]=11'b11101110111;
		Table[239]=11'b11101111111;
		Table[240]=11'b11110000111;
		Table[241]=11'b11110001111;
		Table[242]=11'b11110010111;
		Table[243]=11'b11110011111;
		Table[244]=11'b11110100111;
		Table[245]=11'b11110101111;
		Table[246]=11'b11110110111;
		Table[247]=11'b11110111111;
		Table[248]=11'b11111000111;
		Table[249]=11'b11111001111;
		Table[250]=11'b11111010111;
		Table[251]=11'b11111011111;
		Table[252]=11'b11111100111;
		Table[253]=11'b11111101111;
		Table[254]=11'b11111110111;
		Table[255]=11'b11111111111;
	end
	
	always @(U) begin
		F = Table[U][10:3];
		P = Table[U][2:0];
	end

endmodule
